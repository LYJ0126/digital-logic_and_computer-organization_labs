`timescale 1ns / 1ps


module cache_tb();


//add your code here
endmodule
