module cache_top 
(
    input         rst, 
    input         clk,

    //------gpio-------
    output     [15:0] led,
    input      [15 :0] switch,       
    output reg [7 :0] AN,
    output reg [6 :0] SEG
);

// Add your code here
endmodule
