`timescale 1ns / 1ps

module ALU32(
   output  [31:0] result,      //32λ������
   output  zero,               //���Ϊ0��־λ
   input   [31:0] dataa,      //32λ�������룬�͵�ALU�˿�A   
   input   [31:0] datab,      //32λ�������룬�͵�ALU�˿�B  
   input   [3:0] aluctr      //4λALU���������ź�
); 
//add your code here
endmodule
